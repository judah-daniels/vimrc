Vim�UnDo� �D�IN��k䠪������|����X9J   a          Y                          b�*,    _�                     Q        ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�)�     �   Q   W   S    �   Q   R   S    5�_�                    R       ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�)�     �   Q   T   X          always @(posedge i_clk)5�_�                    R       ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�)�     �   R   T   Z          �   R   T   Y    5�_�                    S       ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�)�     �   R   T   Z      
    ifdef 5�_�                    S       ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�)�     �   R   T   Z      `ifdef 5�_�      
             X   	    ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�*    �   X   Z   [          �   X   Z   Z    5�_�         	       
   Y       ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�*    �   X   Z   [      `enddef5�_�   
                  S        ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�*+    �   S   Z   [    �   S   T   [    5�_�             
   	   Y        ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�*     �   X   Z   [       5�_�              	      Y       ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�*     �   X   Z   [      `endef5�_�                    X   	    ����                                                                                                                                                                                                                                                                                                                            P           N   *       v   d    b�)�     �   X   Y   Z          �   X   Z   [      `endmodule-1-15��
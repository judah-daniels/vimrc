Vim�UnDo� 3�t�Z2y����R?�I!&, M�Ab3ϵ�v   e       always @(posedge i_clk)   ^                          b�    _�                     \       ����                                                                                                                                                                                                                                                                                                                                                             b��'     �   \   ^   f          �   \   ^   e    5�_�                    ]       ����                                                                                                                                                                                                                                                                                                                                                             b��6     �   \   ^   f              else if (i_ce)5�_�                    ]       ����                                                                                                                                                                                                                                                                                                                                                             b��7     �   \   _   f              else if (!i_ce)5�_�                    ]       ����                                                                                                                                                                                                                                                                                                                                                             b��M     �   \   ]                  else if (!i_ce)5�_�                    ]       ����                                                                                                                                                                                                                                                                                                                                                             b��M    �   \   ]                      assert(o_data 5�_�                   Y       ����                                                                                                                                                                                                                                                                                                                                                             b��     �   X   Z   e      "        if (!i_ce && f_past_valid)5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             b��    �   X   Z   e      (        if (!$past(i_ce && f_past_valid)5�_�                    \       ����                                                                                                                                                                                                                                                                                                                                                             b�b     �   \   ^   f          �   \   ^   e    5�_�                    ]       ����                                                                                                                                                                                                                                                                                                                                                             b�i     �   \   ]                  else 5�_�                    ^       ����                                                                                                                                                                                                                                                                                                                                                             b�     �   ]   _   e          always @(posedge i_clk)5�_�                    ^       ����                                                                                                                                                                                                                                                                                                                                                             b�     �   ]   _   e          always @( i_clk)5�_�                     ^       ����                                                                                                                                                                                                                                                                                                                                                             b�    �   ]   _   e          always @( _clk)5�_�                   ]        ����                                                                                                                                                                                                                                                                                                                                                             b��N     �   \   ^   e       5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e      !        if (i_ce && f_past_valid)5�_�      	              Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e               if (_ce && f_past_valid)5�_�      
           	   Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e              if (ce && f_past_valid)5�_�   	              
   Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e              if (e && f_past_valid)5�_�   
                 Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e              if ( && f_past_valid)5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e              if (&& f_past_valid)5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e              if (& f_past_valid)5�_�                    Y       ����                                                                                                                                                                                                                                                                                                                                                             b���     �   X   Z   e              if ( f_past_valid)5�_�                     Y       ����                                                                                                                                                                                                                                                                                                                                                             b���    �   X   Z   e              if (f_past_valid)5��
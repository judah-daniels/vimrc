Vim�UnDo� r&�he�v ���aDy�6e��,4��P X7m   ]           assume(i_reset == 0);   P         %       %   %   %    b�,�    _�                     F       ����                                                                                                                                                                                                                                                                                                                               J          K       v   [    b�*R     �   F   U   O    �   F   G   O    5�_�      	              \        ����                                                                                                                                                                                                                                                                                                                            ]           ]                   b�*a     �   [   \          `endif5�_�      
          	   W        ����                                                                                                                                                                                                                                                                                                                            W           Z           V        b�*�     �   V   W          	always @(*)   		assert(!o_bit);       always @(posedge i_clk)   !        assume(fib_bit==gal_bit);5�_�   	              
   S        ����                                                                                                                                                                                                                                                                                                                            W           W           V        b�*�     �   S   X   X    �   S   T   X    5�_�   
                 Z        ����                                                                                                                                                                                                                                                                                                                            [           [           V        b�*�    �   Y   Z          `ifdef	FORMAL5�_�                    X        ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�*�     �   W   Z   [      `endif5�_�                    Z        ����                                                                                                                                                                                                                                                                                                                            [           [           V        b�*�     �   Y   Z           5�_�                    Q       ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�*�     �   P   R   [      *            assert(o_data == $past(o_data)5�_�                    Q   $    ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�*�     �   P   R   [      +            assert(fib_bit == $past(o_data)5�_�                    R       ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�+$     �   Q   S   [      *                && a_data == $past(a_data)5�_�                    R   !    ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�+'     �   Q   S   [      (                && i_in == $past(a_data)5�_�                    S   #    ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�+(     �   R   T   [      ,                && b_data == $past(b_data));5�_�                    S       ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�+,    �   R   T   [      *                && b_data == $past(i_in));5�_�                    R       ����                                                                                                                                                                                                                                                                                                                            Z           Z           V        b�+7    �   Q   R          &                && i_in == $past(i_in)5�_�                    Q   +    ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�+C    �   P   R   Z      +            assert(fib_bit == $past(fib_bit5�_�                    R   !    ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�+�     �   Q   S   Z      (                && i_in == $past(i_in));5�_�                    R       ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�+�    �   Q   S   Z      +                && i_in == $past(gal_bit));5�_�                    P   (    ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�+�     �   O   Q   Z      )        if (!$past(i_ce) && f_past_valid)5�_�                    P   -    ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�+�    �   O   Q   Z      ;        if (!$past(i_ce) && f_past_valid && !past(i_reset))5�_�                    V       ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�,    �   U   W   Z      !        assume(fib_bit==gal_bit);5�_�                   U       ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�,P    �   T   V   Z          always @(posedge i_clk)5�_�                    M       ����                                                                                                                                                                                                                                                                                                                            Y           Y           V        b�,j     �   M   Q   [          �   M   O   Z    5�_�                    P       ����                                                                                                                                                                                                                                                                                                                            \           \           V        b�,w     �   O   P              -15�_�                     O       ����                                                                                                                                                                                                                                                                                                                            [           [           V        b�,y     �   N   P   \          assume @(*)5�_�      "               O   	    ����                                                                                                                                                                                                                                                                                                                            [           [           V        b�,|     �   O   Q   ]              �   O   Q   \    5�_�       #   !       "   P       ����                                                                                                                                                                                                                                                                                                                            \           \           V        b�,�     �   O   Q   ]              assumme(i_reset == 0);5�_�   "   $           #   P       ����                                                                                                                                                                                                                                                                                                                            \           \           V        b�,�     �   P   R   ^          �   P   R   ]    5�_�   #   %           $   Q       ����                                                                                                                                                                                                                                                                                                                            ]           ]           V        b�,�     �   P   Q              -15�_�   $               %   P       ����                                                                                                                                                                                                                                                                                                                            \           \           V        b�,�    �   O   Q   ]              assume(i_reset == 0);5�_�               "   !   P       ����                                                                                                                                                                                                                                                                                                                            \           \           V        b�,�     �   O   Q   ]              assmme(i_reset == 0);5�_�                    U       ����                                                                                                                                                                                                                                                                                                                            X           X           V        b�,<   
 �   T   V        5�_�            	      V        ����                                                                                                                                                                                                                                                                                                                            Z           V                   b�*{     �   U   [   \      ifdef	FORMAL      always @(*)      	assert(!o_bit);      always @(posedge i_clk)           assume(fib_bit==gal_bit);5�_�                    V        ����                                                                                                                                                                                                                                                                                                                            X           V                   b�*}     �   U   X        5�_�                    V       ����                                                                                                                                                                                                                                                                                                                            W           V                   b�*~     �   U   W        5�_�                    V       ����                                                                                                                                                                                                                                                                                                                            V           V                   b�*~     �   U   W        5�_�                     V       ����                                                                                                                                                                                                                                                                                                                            V           V                   b�*    �   U   W        5�_�                    U        ����                                                                                                                                                                                                                                                                                                                            [           U                   b�*h     �   T   \   \          ifdef	FORMAL      always @(*)      	assert(!o_bit);      always @(posedge i_clk)           assume(fib_bit==gal_bit);    5��